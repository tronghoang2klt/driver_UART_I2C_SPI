library ieee;
use	ieee.std_logic_1164.all;
library std;
use	std.standard.all;
library work;
use 	work.all;
entity Slave_SPI is
port(
	i_clk	: in std_logic
	----------MOSI------
	----------MISO------
	----------4 wire----
	
);
end Slave_SPI;
architecture main of Slave_SPI is
begin
end main;